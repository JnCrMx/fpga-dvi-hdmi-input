module tmds_decoder (
  input logic [9:0] tmds_symbol,

  output logic valid,
  output logic [7:0] channel_data,
  output logic [1:0] c,
  output logic de
);

logic [9:0] tmp_tmds_symbol;

always_comb begin
  c = 0;
  channel_data = 0;
  tmp_tmds_symbol = 0;
  de = 0; // assume control
  valid = 0;

  case (tmds_symbol[9:0])
    10'b1101010100: c = 2'b00;
    10'b0010101011: c = 2'b01;
    10'b0101010100: c = 2'b10;
    10'b1010101011: c = 2'b11;
    default: begin
      de = 1; // and if it is not control, then it is data
      if (tmds_symbol[9] == 1) begin
        tmp_tmds_symbol = {tmds_symbol[9:8], ~tmds_symbol[7:0]};
      end else begin
        tmp_tmds_symbol = tmds_symbol;
      end
      if (tmds_symbol[8] == 1) begin
        channel_data[0] = tmp_tmds_symbol[0];
        channel_data[1] = tmp_tmds_symbol[1] ^ tmp_tmds_symbol[0];
        channel_data[2] = tmp_tmds_symbol[2] ^ tmp_tmds_symbol[1];
        channel_data[3] = tmp_tmds_symbol[3] ^ tmp_tmds_symbol[2];
        channel_data[4] = tmp_tmds_symbol[4] ^ tmp_tmds_symbol[3];
        channel_data[5] = tmp_tmds_symbol[5] ^ tmp_tmds_symbol[4];
        channel_data[6] = tmp_tmds_symbol[6] ^ tmp_tmds_symbol[5];
        channel_data[7] = tmp_tmds_symbol[7] ^ tmp_tmds_symbol[6];
      end else begin
        channel_data[0] = tmp_tmds_symbol[0];
        channel_data[1] = ~(tmp_tmds_symbol[1] ^ tmp_tmds_symbol[0]);
        channel_data[2] = ~(tmp_tmds_symbol[2] ^ tmp_tmds_symbol[1]);
        channel_data[3] = ~(tmp_tmds_symbol[3] ^ tmp_tmds_symbol[2]);
        channel_data[4] = ~(tmp_tmds_symbol[4] ^ tmp_tmds_symbol[3]);
        channel_data[5] = ~(tmp_tmds_symbol[5] ^ tmp_tmds_symbol[4]);
        channel_data[6] = ~(tmp_tmds_symbol[6] ^ tmp_tmds_symbol[5]);
        channel_data[7] = ~(tmp_tmds_symbol[7] ^ tmp_tmds_symbol[6]);
      end
    end
  endcase

  //valid (Data values generated by python script)
  case (tmds_symbol)
    `include "../../../build/tmds_valid/generate/fragments/valid_tmds.sv"

    //Ctrl
    10'b0010101011: valid = 1;
    10'b0101010100: valid = 1;
    10'b1010101011: valid = 1;
    10'b1101010100: valid = 1;

    default: valid = 0;
  endcase
end

endmodule
